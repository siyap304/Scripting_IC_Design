`timescale 1ns / 1ps
module LAB1_using_decoder(
    input [4:0] A,
    output OUT,
    input [2:0] S);

    wire [31:0] I;
    wire [9:2] M;
    wire [31:0] X;
    
    or(M[2], ~S[2], S[1], ~S[0]);
    or(M[3], ~S[2], S[1], S[0]);
    or(M[4], S[2], ~S[1], ~S[0]);
    or(M[5], S[2], ~S[1], S[0]);
    or(M[6], S[2], S[1], ~S[0]);
    or(M[7], S[2], S[1], S[0]);
    or(M[8], ~S[2], ~S[1], ~S[0]);
    or(M[9], ~S[2], ~S[1], S[0]);
    
    assign X = 32'b0;
    assign I = 32'b0;
    
    or(X[0], M[2], M[3], M[4], M[5], M[6], M[7], M[8], M[9]);
    or(X[2], M[2]);
    or(X[3], M[3]);
    or(X[4], M[2], M[4]);
    or(X[5], M[5]);
    or(X[6], M[2], M[3], M[6]);
    or(X[7], M[7]);
    or(X[8], M[2], M[4], M[8]);
    or(X[9], M[9]);
    or(X[10], M[2], M[5]);
    or(X[12], M[2], M[4], M[3], M[6]);
    or(X[14], M[2], M[7]);
    or(X[15], M[3], M[5]);
    or(X[16], M[2], M[4], M[8]);
    or(X[18], M[2], M[3], M[6], M[9]);
    or(X[20], M[2], M[4], M[5]);
    or(X[21], M[3], M[7]);
    or(X[22], M[2]);
    or(X[24], M[2], M[3], M[4], M[6], M[8]);
    or(X[25], M[5]);
    or(X[26], M[2]);
    or(X[27], M[3], M[9]);
    or(X[28], M[2], M[4], M[7]);
    or(X[30], M[2], M[3], M[5], M[6]);
    
    and(I[0], ~A[4], ~A[3], ~A[2], ~A[1], ~A[0], X[0]);
    and(I[2], ~A[4], ~A[3], ~A[2], A[1], ~A[0], X[2]);
    and(I[3], ~A[4], ~A[3], ~A[2], A[1], A[0], X[3]);
    and(I[4], ~A[4], ~A[3], A[2], ~A[1], ~A[0], X[4]);
    and(I[5], ~A[4], ~A[3], A[2], ~A[1], A[0], X[5]);
    and(I[6], ~A[4], ~A[3], A[2], A[1], ~A[0], X[6]);
    and(I[7], ~A[4], ~A[3], A[2], A[1], A[0], X[7]);
    and(I[8], ~A[4], A[3], ~A[2], ~A[1], ~A[0], X[8]);
    and(I[9], ~A[4], A[3], ~A[2], ~A[1], A[0], X[9]);
    and(I[10], ~A[4], A[3], ~A[2], A[1], ~A[0], X[10]);
    and(I[12], ~A[4], A[3], A[2], ~A[1], ~A[0], X[12]);
    and(I[14], ~A[4], A[3], A[2], A[1], ~A[0], X[14]);
    and(I[15], ~A[4], A[3], A[2], A[1], A[0], X[15]);
    and(I[16], A[4], ~A[3], ~A[2], ~A[1], ~A[0], X[16]);
    and(I[18], A[4], ~A[3], ~A[2], A[1], ~A[0], X[18]);
    and(I[20], A[4], ~A[3], A[2], ~A[1], ~A[0], X[20]);
    and(I[21], A[4], ~A[3], A[2], ~A[1], A[0], X[21]);
    and(I[22], A[4], ~A[3], A[2], A[1], ~A[0], X[22]);
    and(I[24], A[4], A[3], ~A[2], ~A[1], ~A[0], X[24]);
    and(I[25], A[4], A[3], ~A[2], ~A[1], A[0], X[25]);
    and(I[26], A[4], A[3], ~A[2], A[1], ~A[0], X[26]);
    and(I[27], A[4], A[3], ~A[2], A[1], A[0], X[27]);
    and(I[28], A[4], A[3], A[2], ~A[1], ~A[0], X[28]);
    and(I[30], A[4], A[3], A[2], A[1], ~A[0], X[30]);
    
endmodule
